module top_module (
    input [2:0] a,
    output [15:0] q ); 
    // m1 + m6
    assign q[15] = (~a[2] & ~a[1] & a[0]) | (a[2] & a[1] & ~a[0]);
    // m3 + m5 + m6
    assign q[14] = (~a[2] & a[1] & a[0]) | (a[2] & ~a[1] & a[0]) | (a[2] & a[1] & ~a[0]);
    // m1 + m2 + (m4 + m5) + m7
    assign q[13] = (~a[2] & ~a[1] & a[0]) | (~a[2] & a[1] & ~a[0]) | (a[2] & ~a[1]) | (a[2] & a[1] & a[0]);
    // m0 + m3 
    assign q[12] = ~a[2] & (a[1] ~^ a[0]);
    // m1 + m3 + m7
    assign q[11] = (~a[2] & a[0]) | (a[1] & a[0]);
    // (m1 + m5) | (m2 + m6) | m7
    assign q[10] = (~a[1] & a[0]) | (a[1] & ~a[0]) | (a[2] & a[1] & a[0]);
    // (m0 + m1 + m2 + m3) + m7
    assign q[9] = ~a[2] | (a[1] & a[0]);
    // (m6 + m7) + (m2 + m6)
    assign q[8] = (a[2] & a[1]) | (a[1] & ~a[0]);
    // (m1 + m5) + m2
    assign q[7] = (~a[1] & a[0]) | (~a[2] & a[1] & ~a[0]);
    //(m1 + m5) + (m4 + m5) + m2
    assign q[6] = (~a[1] & a[0]) | (a[2] & ~a[1]) | (~a[2] & a[1] & ~a[0]);
    // (m0 + m1) + (m4 + m6)
    assign q[5] = (~a[2] & ~a[1]) | (a[2] & ~a[0]);
    // m0 + m7 + m2
    assign q[4] = (~a[2] & ~a[1] & ~a[0]) | (a[2] & a[1] & a[0]) | (~a[2] & a[1] & ~a[0]);
    // (m3 + m5) + (m3 + m7)
    assign q[3] = (a[2] & a[0]) | (a[1] & a[0]);
    // (m2 + m3 + m4 + m5) + (m5 + m6)
    assign q[2] = (a[2] ^ a[1]) | (a[2] & ~a[0]);
    // (m0 + m4) | (m4 + m6) | (m3 + m5)
    assign q[1] = (~a[1] & ~a[0]) | (a[2] & ~a[0]) | ((a[2] ^ a[1]) & a[0]);
    // m7
    assign q[0] = (a[2] & a[1] & a[0]);
endmodule